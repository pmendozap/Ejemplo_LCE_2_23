.TITLE Circuito ohm
.OP
V1 N1 0 10
R1 N1 0 1k
.END